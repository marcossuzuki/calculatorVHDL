library verilog;
use verilog.vl_types.all;
entity somador_for_vlg_vec_tst is
end somador_for_vlg_vec_tst;
