library verilog;
use verilog.vl_types.all;
entity PWM_vlg_vec_tst is
end PWM_vlg_vec_tst;
