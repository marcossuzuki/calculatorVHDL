library verilog;
use verilog.vl_types.all;
entity clock_div_vlg_vec_tst is
end clock_div_vlg_vec_tst;
